`define MD_OP_MUL 1'b0
`define MD_OP_DIV 1'b1

`define MD_OUT_LO  1'b0
`define MD_OUT_HI  1'b1

